`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2015/07/09 14:26:01
// Design Name: 
// Module Name: PIC16F54
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PIC16F54(

    );
    
    
    ALU8    ALU8_01(
    );
    
    Reg_File    Reg_File_01(
    );
endmodule
